// `default_nettype none
// `include "def.sv"

// module alu


// endmodule

// `default_nettype wire
