// `default_nettype none
// `include "def.sv"

// module fetch



// endmodule

// `default_nettype wire
